module top ();

design_1 design_1_wrapper
   (
    clk_200(),
    sys_arstn(),
    S_AXIS_1_tdata(),
    S_AXIS_1_tlast(),
    S_AXIS_1_tready(),
    S_AXIS_1_tvalid()
    );

endmodule